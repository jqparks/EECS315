*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'jqp' on Thu Feb 25 2016 at 10:06:25

*
* Globals.
*
.global GND VDD

*
* MAIN CELL: Component pathname : /home/jqp/eecs315/lab2/dff
*
        MP12 BCLK BCLK- VDD VDD p L=2u W=18u
        MP11 BCLK- CLK VDD VDD p L=2u W=18u
        MN15 QB N$62 GND GND n L=2u W=10u
        MP4 N$10 D VDD VDD p L=2u W=27u
        MN12 BCLK BCLK- GND GND n L=2u W=10u
        MN11 BCLK- CLK GND GND n L=2u W=10u
        MN10 N$101 N$62 GND GND n L=2u W=5u
        MN9 N$68 N$101 GND GND n L=2u W=5u
        MN8 N$62 BCLK- N$68 GND n L=2u W=5u
        MN7 N$66 N$26 GND GND n L=2u W=15u
        MN6 N$62 BCLK N$66 GND n L=2u W=15u
        MN5 N$31 N$26 GND GND n L=2u W=5u
        MN4 N$54 N$31 GND GND n L=2u W=5u
        MN3 N$56 D GND GND n L=2u W=15u
        MN2 N$26 BCLK N$54 GND n L=2u W=5u
        MN1 N$26 BCLK- N$56 GND n L=2u W=15u
        MP10 N$101 N$62 VDD VDD p L=2u W=5u
        MP9 N$62 BCLK N$24 VDD p L=2u W=5u
        MP8 N$62 BCLK- N$22 VDD p L=2u W=27u
        MP7 N$24 N$101 VDD VDD p L=2u W=5u
        MP6 N$22 N$26 VDD VDD p L=2u W=27u
        MP5 N$12 N$31 VDD VDD p L=2u W=5u
        MN16 Q QB GND GND n L=2u W=10u
        MP3 N$26 BCLK N$10 VDD p L=2u W=27u
        MP2 N$31 N$26 VDD VDD p L=2u W=5u
        MP1 N$26 BCLK- N$12 VDD p L=2u W=5u
        MP14 Q QB VDD VDD p L=2u W=18u
        MP13 QB N$62 VDD VDD p L=2u W=18u
*
.end

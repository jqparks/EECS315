*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'jqp' on Wed Feb 24 2016 at 11:44:13

*
* Globals.
*
.global GND VDD

*
* MAIN CELL: Component pathname : /home/jqp/eecs315/lab2/aoi
*
        MN4 N$28 B1 GND GND n L=2u W=10u
        MN3 N$26 A1 GND GND n L=2u W=10u
        MN2 OUTPUT B0 N$28 GND n L=2u W=10u
        MN1 OUTPUT A0 N$26 GND n L=2u W=10u
        MP2 OUTPUT B1 N$18 VDD p L=2u W=13u
        MP4 N$18 A1 VDD VDD p L=2u W=13u
        MP3 N$18 A0 VDD VDD p L=2u W=13u
        MP1 OUTPUT B0 N$18 VDD p L=2u W=13u
*
.end

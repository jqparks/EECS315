* Component: /home/jqp/eecs315/lab2/aoi  Viewpoint: ami05a
.INCLUDE /home/jqp/eecs315/lab2/aoi/ami05a/aoi_ami05a.spi
.LIB /mgc/adk3_1/technology/ic/models/VDD_5.mod
.LIB /mgc/adk3_1/technology/ic/models/ami05.mod
.PROBE TRAN V(A0) V(A1) V(B0) V(B1)
.PROBE TRAN V(OUTPUT)

VFORCE__A0 A0 GND pulse (0 5 0 1e-09 1e-09 25n 50n)

VFORCE__A1 A1 GND pulse (0 5 0 1e-09 1e-09 50n 100n)

VFORCE__B0 B0 GND pulse (0 5 0 1e-09 1e-09 100n 200n)

VFORCE__B1 B1 GND pulse (0 5 0 1e-09 1e-09 200n 400n)




.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

.TEMP 27 

.TRAN  0 800n 0n 

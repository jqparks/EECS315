*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'jqp' on Mon Feb 22 2016 at 21:40:23

*
* Globals.
*
.global GND VDD

*
* MAIN CELL: Component pathname : /home/jqp/eecs315/lab2/nand
*
        MN2 N$5 INPUT2 GND GND n L=2u W=10u
        MN1 OUTPUT INPUT1 N$5 GND n L=2u W=10u
        MP2 OUTPUT INPUT2 VDD VDD p L=2u W=12u
        MP1 OUTPUT INPUT1 VDD VDD p L=2u W=12u
*
.end
